magic
tech gf180mcuC
magscale 1 5
timestamp 1670256780
<< obsm1 >>
rect 672 1538 29895 28321
<< metal2 >>
rect 980 29600 1092 29900
rect 1988 29600 2100 29900
rect 2996 29600 3108 29900
rect 4004 29600 4116 29900
rect 5012 29600 5124 29900
rect 6020 29600 6132 29900
rect 7028 29600 7140 29900
rect 8036 29600 8148 29900
rect 9044 29600 9156 29900
rect 10388 29600 10500 29900
rect 11396 29600 11508 29900
rect 12404 29600 12516 29900
rect 13412 29600 13524 29900
rect 14420 29600 14532 29900
rect 15428 29600 15540 29900
rect 16436 29600 16548 29900
rect 17444 29600 17556 29900
rect 18452 29600 18564 29900
rect 19460 29600 19572 29900
rect 20804 29600 20916 29900
rect 21812 29600 21924 29900
rect 22820 29600 22932 29900
rect 23828 29600 23940 29900
rect 24836 29600 24948 29900
rect 25844 29600 25956 29900
rect 26852 29600 26964 29900
rect 27860 29600 27972 29900
rect 28868 29600 28980 29900
rect 29876 29600 29988 29900
rect -28 100 84 400
rect 980 100 1092 400
rect 1988 100 2100 400
rect 2996 100 3108 400
rect 4004 100 4116 400
rect 5012 100 5124 400
rect 6020 100 6132 400
rect 7028 100 7140 400
rect 8036 100 8148 400
rect 9044 100 9156 400
rect 10388 100 10500 400
rect 11396 100 11508 400
rect 12404 100 12516 400
rect 13412 100 13524 400
rect 14420 100 14532 400
rect 15428 100 15540 400
rect 16436 100 16548 400
rect 17444 100 17556 400
rect 18452 100 18564 400
rect 19460 100 19572 400
rect 20804 100 20916 400
rect 21812 100 21924 400
rect 22820 100 22932 400
rect 23828 100 23940 400
rect 24836 100 24948 400
rect 25844 100 25956 400
rect 26852 100 26964 400
rect 27860 100 27972 400
rect 28868 100 28980 400
<< obsm2 >>
rect 70 29930 29890 29951
rect 70 29570 950 29930
rect 1122 29570 1958 29930
rect 2130 29570 2966 29930
rect 3138 29570 3974 29930
rect 4146 29570 4982 29930
rect 5154 29570 5990 29930
rect 6162 29570 6998 29930
rect 7170 29570 8006 29930
rect 8178 29570 9014 29930
rect 9186 29570 10358 29930
rect 10530 29570 11366 29930
rect 11538 29570 12374 29930
rect 12546 29570 13382 29930
rect 13554 29570 14390 29930
rect 14562 29570 15398 29930
rect 15570 29570 16406 29930
rect 16578 29570 17414 29930
rect 17586 29570 18422 29930
rect 18594 29570 19430 29930
rect 19602 29570 20774 29930
rect 20946 29570 21782 29930
rect 21954 29570 22790 29930
rect 22962 29570 23798 29930
rect 23970 29570 24806 29930
rect 24978 29570 25814 29930
rect 25986 29570 26822 29930
rect 26994 29570 27830 29930
rect 28002 29570 28838 29930
rect 29010 29570 29846 29930
rect 70 430 29890 29570
rect 114 350 950 430
rect 1122 350 1958 430
rect 2130 350 2966 430
rect 3138 350 3974 430
rect 4146 350 4982 430
rect 5154 350 5990 430
rect 6162 350 6998 430
rect 7170 350 8006 430
rect 8178 350 9014 430
rect 9186 350 10358 430
rect 10530 350 11366 430
rect 11538 350 12374 430
rect 12546 350 13382 430
rect 13554 350 14390 430
rect 14562 350 15398 430
rect 15570 350 16406 430
rect 16578 350 17414 430
rect 17586 350 18422 430
rect 18594 350 19430 430
rect 19602 350 20774 430
rect 20946 350 21782 430
rect 21954 350 22790 430
rect 22962 350 23798 430
rect 23970 350 24806 430
rect 24978 350 25814 430
rect 25986 350 26822 430
rect 26994 350 27830 430
rect 28002 350 28838 430
rect 29010 350 29890 430
<< metal3 >>
rect 100 29876 400 29988
rect 100 28868 400 28980
rect 29600 28868 29900 28980
rect 100 27860 400 27972
rect 29600 27860 29900 27972
rect 100 26852 400 26964
rect 29600 26852 29900 26964
rect 100 25844 400 25956
rect 29600 25844 29900 25956
rect 100 24836 400 24948
rect 29600 24836 29900 24948
rect 100 23828 400 23940
rect 29600 23828 29900 23940
rect 100 22820 400 22932
rect 29600 22820 29900 22932
rect 100 21812 400 21924
rect 29600 21812 29900 21924
rect 100 20804 400 20916
rect 29600 20804 29900 20916
rect 100 19460 400 19572
rect 29600 19460 29900 19572
rect 100 18452 400 18564
rect 29600 18452 29900 18564
rect 100 17444 400 17556
rect 29600 17444 29900 17556
rect 100 16436 400 16548
rect 29600 16436 29900 16548
rect 100 15428 400 15540
rect 29600 15428 29900 15540
rect 100 14420 400 14532
rect 29600 14420 29900 14532
rect 100 13412 400 13524
rect 29600 13412 29900 13524
rect 100 12404 400 12516
rect 29600 12404 29900 12516
rect 100 11396 400 11508
rect 29600 11396 29900 11508
rect 100 10388 400 10500
rect 29600 10388 29900 10500
rect 100 9044 400 9156
rect 29600 9044 29900 9156
rect 100 8036 400 8148
rect 29600 8036 29900 8148
rect 100 7028 400 7140
rect 29600 7028 29900 7140
rect 100 6020 400 6132
rect 29600 6020 29900 6132
rect 100 5012 400 5124
rect 29600 5012 29900 5124
rect 100 4004 400 4116
rect 29600 4004 29900 4116
rect 100 2996 400 3108
rect 29600 2996 29900 3108
rect 100 1988 400 2100
rect 29600 1988 29900 2100
rect 100 980 400 1092
rect 29600 980 29900 1092
rect 29600 -28 29900 84
<< obsm3 >>
rect 430 29846 29666 29946
rect 350 29010 29666 29846
rect 430 28838 29570 29010
rect 350 28002 29666 28838
rect 430 27830 29570 28002
rect 350 26994 29666 27830
rect 430 26822 29570 26994
rect 350 25986 29666 26822
rect 430 25814 29570 25986
rect 350 24978 29666 25814
rect 430 24806 29570 24978
rect 350 23970 29666 24806
rect 430 23798 29570 23970
rect 350 22962 29666 23798
rect 430 22790 29570 22962
rect 350 21954 29666 22790
rect 430 21782 29570 21954
rect 350 20946 29666 21782
rect 430 20774 29570 20946
rect 350 19602 29666 20774
rect 430 19430 29570 19602
rect 350 18594 29666 19430
rect 430 18422 29570 18594
rect 350 17586 29666 18422
rect 430 17414 29570 17586
rect 350 16578 29666 17414
rect 430 16406 29570 16578
rect 350 15570 29666 16406
rect 430 15398 29570 15570
rect 350 14562 29666 15398
rect 430 14390 29570 14562
rect 350 13554 29666 14390
rect 430 13382 29570 13554
rect 350 12546 29666 13382
rect 430 12374 29570 12546
rect 350 11538 29666 12374
rect 430 11366 29570 11538
rect 350 10530 29666 11366
rect 430 10358 29570 10530
rect 350 9186 29666 10358
rect 430 9014 29570 9186
rect 350 8178 29666 9014
rect 430 8006 29570 8178
rect 350 7170 29666 8006
rect 430 6998 29570 7170
rect 350 6162 29666 6998
rect 430 5990 29570 6162
rect 350 5154 29666 5990
rect 430 4982 29570 5154
rect 350 4146 29666 4982
rect 430 3974 29570 4146
rect 350 3138 29666 3974
rect 430 2966 29570 3138
rect 350 2130 29666 2966
rect 430 1958 29570 2130
rect 350 1122 29666 1958
rect 430 950 29570 1122
rect 350 114 29666 950
rect 350 70 29570 114
<< metal4 >>
rect 2224 1538 2384 28254
rect 9904 1538 10064 28254
rect 17584 1538 17744 28254
rect 25264 1538 25424 28254
<< labels >>
rlabel metal3 s 29600 28868 29900 28980 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 29600 7028 29900 7140 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 2996 29600 3108 29900 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 100 16436 400 16548 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 26852 29600 26964 29900 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 21812 29600 21924 29900 6 io_in[14]
port 6 nsew signal input
rlabel metal3 s 100 18452 400 18564 6 io_in[15]
port 7 nsew signal input
rlabel metal3 s 100 5012 400 5124 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 10388 29600 10500 29900 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 8036 100 8148 400 6 io_in[18]
port 10 nsew signal input
rlabel metal3 s 100 4004 400 4116 6 io_in[19]
port 11 nsew signal input
rlabel metal3 s 29600 26852 29900 26964 6 io_in[1]
port 12 nsew signal input
rlabel metal3 s 29600 980 29900 1092 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 25844 29600 25956 29900 6 io_in[21]
port 14 nsew signal input
rlabel metal3 s 100 20804 400 20916 6 io_in[22]
port 15 nsew signal input
rlabel metal3 s 100 26852 400 26964 6 io_in[23]
port 16 nsew signal input
rlabel metal3 s 29600 13412 29900 13524 6 io_in[24]
port 17 nsew signal input
rlabel metal3 s 100 2996 400 3108 6 io_in[25]
port 18 nsew signal input
rlabel metal3 s 100 27860 400 27972 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 14420 29600 14532 29900 6 io_in[27]
port 20 nsew signal input
rlabel metal3 s 29600 27860 29900 27972 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 28868 100 28980 400 6 io_in[29]
port 22 nsew signal input
rlabel metal3 s 29600 9044 29900 9156 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 13412 29600 13524 29900 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 18452 100 18564 400 6 io_in[31]
port 25 nsew signal input
rlabel metal3 s 29600 15428 29900 15540 6 io_in[32]
port 26 nsew signal input
rlabel metal3 s 100 17444 400 17556 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 7028 100 7140 400 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 11396 100 11508 400 6 io_in[35]
port 29 nsew signal input
rlabel metal3 s 29600 2996 29900 3108 6 io_in[36]
port 30 nsew signal input
rlabel metal3 s 100 22820 400 22932 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 9044 29600 9156 29900 6 io_in[3]
port 32 nsew signal input
rlabel metal3 s 29600 10388 29900 10500 6 io_in[4]
port 33 nsew signal input
rlabel metal3 s 29600 16436 29900 16548 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 16436 29600 16548 29900 6 io_in[6]
port 35 nsew signal input
rlabel metal3 s 29600 12404 29900 12516 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 17444 29600 17556 29900 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 19460 29600 19572 29900 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 23828 29600 23940 29900 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 29876 29600 29988 29900 6 io_oeb[10]
port 40 nsew signal output
rlabel metal3 s 29600 24836 29900 24948 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 4004 100 4116 400 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 5012 29600 5124 29900 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 13412 100 13524 400 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 17444 100 17556 400 6 io_oeb[15]
port 45 nsew signal output
rlabel metal3 s 29600 25844 29900 25956 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 26852 100 26964 400 6 io_oeb[17]
port 47 nsew signal output
rlabel metal3 s 29600 19460 29900 19572 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 12404 29600 12516 29900 6 io_oeb[19]
port 49 nsew signal output
rlabel metal3 s 100 14420 400 14532 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 7028 29600 7140 29900 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 15428 29600 15540 29900 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 23828 100 23940 400 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 9044 100 9156 400 6 io_oeb[23]
port 54 nsew signal output
rlabel metal3 s 29600 8036 29900 8148 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 8036 29600 8148 29900 6 io_oeb[25]
port 56 nsew signal output
rlabel metal3 s 29600 20804 29900 20916 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 1988 100 2100 400 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 27860 100 27972 400 6 io_oeb[28]
port 59 nsew signal output
rlabel metal3 s 29600 6020 29900 6132 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 28868 29600 28980 29900 6 io_oeb[2]
port 61 nsew signal output
rlabel metal3 s 100 24836 400 24948 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 24836 100 24948 400 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 12404 100 12516 400 6 io_oeb[32]
port 64 nsew signal output
rlabel metal3 s 100 23828 400 23940 6 io_oeb[33]
port 65 nsew signal output
rlabel metal3 s 29600 22820 29900 22932 6 io_oeb[34]
port 66 nsew signal output
rlabel metal3 s 100 13412 400 13524 6 io_oeb[35]
port 67 nsew signal output
rlabel metal3 s 29600 1988 29900 2100 6 io_oeb[36]
port 68 nsew signal output
rlabel metal3 s 100 29876 400 29988 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 4004 29600 4116 29900 6 io_oeb[3]
port 70 nsew signal output
rlabel metal3 s 100 19460 400 19572 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 21812 100 21924 400 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 2996 100 3108 400 6 io_oeb[6]
port 73 nsew signal output
rlabel metal3 s 100 12404 400 12516 6 io_oeb[7]
port 74 nsew signal output
rlabel metal3 s 29600 -28 29900 84 6 io_oeb[8]
port 75 nsew signal output
rlabel metal3 s 29600 17444 29900 17556 6 io_oeb[9]
port 76 nsew signal output
rlabel metal3 s 29600 11396 29900 11508 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 22820 100 22932 400 6 io_out[10]
port 78 nsew signal output
rlabel metal3 s 100 21812 400 21924 6 io_out[11]
port 79 nsew signal output
rlabel metal3 s 29600 5012 29900 5124 6 io_out[12]
port 80 nsew signal output
rlabel metal3 s 100 15428 400 15540 6 io_out[13]
port 81 nsew signal output
rlabel metal3 s 100 980 400 1092 6 io_out[14]
port 82 nsew signal output
rlabel metal3 s 29600 21812 29900 21924 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 25844 100 25956 400 6 io_out[16]
port 84 nsew signal output
rlabel metal3 s 29600 23828 29900 23940 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 15428 100 15540 400 6 io_out[18]
port 86 nsew signal output
rlabel metal3 s 100 6020 400 6132 6 io_out[19]
port 87 nsew signal output
rlabel metal3 s 100 11396 400 11508 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s -28 100 84 400 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 19460 100 19572 400 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 1988 29600 2100 29900 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 11396 29600 11508 29900 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 20804 29600 20916 29900 6 io_out[24]
port 93 nsew signal output
rlabel metal3 s 100 1988 400 2100 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 5012 100 5124 400 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 980 100 1092 400 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 24836 29600 24948 29900 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 18452 29600 18564 29900 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 14420 100 14532 400 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 27860 29600 27972 29900 6 io_out[30]
port 100 nsew signal output
rlabel metal3 s 29600 4004 29900 4116 6 io_out[31]
port 101 nsew signal output
rlabel metal3 s 100 28868 400 28980 6 io_out[32]
port 102 nsew signal output
rlabel metal3 s 100 10388 400 10500 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 6020 100 6132 400 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 10388 100 10500 400 6 io_out[35]
port 105 nsew signal output
rlabel metal3 s 100 9044 400 9156 6 io_out[36]
port 106 nsew signal output
rlabel metal3 s 29600 18452 29900 18564 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 16436 100 16548 400 6 io_out[3]
port 108 nsew signal output
rlabel metal3 s 100 7028 400 7140 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 22820 29600 22932 29900 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 980 29600 1092 29900 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 6020 29600 6132 29900 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 20804 100 20916 400 6 io_out[8]
port 113 nsew signal output
rlabel metal3 s 100 8036 400 8148 6 io_out[9]
port 114 nsew signal output
rlabel metal4 s 2224 1538 2384 28254 6 vdd
port 115 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 28254 6 vdd
port 115 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 28254 6 vss
port 116 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 28254 6 vss
port 116 nsew ground bidirectional
rlabel metal3 s 100 25844 400 25956 6 wb_clk_i
port 117 nsew signal input
rlabel metal3 s 29600 14420 29900 14532 6 wb_rst_i
port 118 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 30000 30000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 421520
string GDS_FILE /home/mm4uz/asic/gf180-shuttle-0/gf180-mul-8-seq/openlane/wrapped_multiplier_8/runs/22_12_05_11_12/results/signoff/wrapped_multiplier_8.magic.gds
string GDS_START 50130
<< end >>

